//7 segment decoder 4bit

module decoder_7segment_4bit(m,out);
	input [3:0] m;
	output [6:0] out;

	assign out = (m==4'b0000) ? (7'b1000000) :
					 (m==4'b0001) ? (7'b1111001) :
					 (m==4'b0010) ? (7'b0100100) :
					 (m==4'b0011) ? (7'b0110000) :
					 (m==4'b0100) ? (7'b0011001) :
					 (m==4'b0101) ? (7'b0010010) :
					 (m==4'b0110) ? (7'b0000010) :
					 (m==4'b0111) ? (7'b1111000) :
					 (m==4'b1000) ? (7'b0000000) :		
					 (m==4'b1001) ? (7'b0010000) :
					 (m==4'b1010) ? (7'b1111111) :
					 (m==4'b1011) ? (7'b1111111) :
					 (m==4'b1100) ? (7'b1111111) :
					 (m==4'b1101) ? (7'b1111111) :
					 (m==4'b1110) ? (7'b1111111) :
					 (m==4'b1111) ? (7'b1111111) :
					 1'bx;
					 
endmodule