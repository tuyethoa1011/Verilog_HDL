library verilog;
use verilog.vl_types.all;
entity morsecode_encoder_vlg_vec_tst is
end morsecode_encoder_vlg_vec_tst;
