library verilog;
use verilog.vl_types.all;
entity morse_code_vlg_vec_tst is
end morse_code_vlg_vec_tst;
