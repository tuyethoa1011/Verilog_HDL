library verilog;
use verilog.vl_types.all;
entity morsecode_shiftregister_vlg_vec_tst is
end morsecode_shiftregister_vlg_vec_tst;
