library verilog;
use verilog.vl_types.all;
entity morsecode_lengthcounter_vlg_vec_tst is
end morsecode_lengthcounter_vlg_vec_tst;
